`ifndef __GLOBALS__
`define __GLOBALS__

// UVM Globals
localparam string IQ_IN_NAME = "../data/read_iq.txt";
localparam string LEFT_OUT_NAME = "../data/left_out_uvm.txt";
localparam string RIGHT_OUT_NAME = "../data/right_out_uvm.txt";
localparam string RIGHT_CMP_NAME = "../data/right_volume.txt";
localparam string LEFT_CMP_NAME = "../data/left_volume.txt";
localparam int CLOCK_PERIOD = 10;

`endif
